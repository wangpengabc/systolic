
module test;
  initial begin
    $display("test!");
    $finish;
  end
endmodule
