
module SubmoduleC(
    input  io_in
);
endmodule
    